/* OR 회로 설계 */
module ORgate(A, B, F);
  input A, B;
  output F;

  assign F=A|B;

endmodule
