/* NOT 회로 설계 */
module NOTgate(A, F);
  input A;
  output F;

  assign F=~A;

endmodule
